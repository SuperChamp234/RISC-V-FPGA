module sev_seg_disp();

endmodule