module RISC_V;

endmodule